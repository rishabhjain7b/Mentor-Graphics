package my_package;

typedef enum{red,green,blue}color;

typedef struct{
	int field_a;
	color c;
	}mystruct;
	
endpackage

