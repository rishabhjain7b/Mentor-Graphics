`define CLK_PERIOD 10
`define REGISTER_WIDTH 32
`define INSTR_WIDTH 32
`define IMMEDIATE_WIDTH 16
`define MEM_READ 3'b101
`define MEM_WRITE 3'b100
`define ARITH_LOGIC 3'b001
`define SHIFT_REG 3'b000

// ARITHMETIC 3'b000
`define 3'b001
ADD 3'b010
`define 3'b011
HADD 3'b100
`define 3'b101
SUB 3'b110
`define 3'b111
NOT 
`define 
AND 
 `define 
OR 
`define 
XOR 
`define 
LHG 
// SHIFTING SHLEFTLOG 3'b000
`define SHLEFTART 3'b001
`define SHRGHTLOG 3'b010
`define SHRGHTART 3'b011
`define 
// DATA TRANSFER 3'b000
`define 3'b100
LOADBYTE 3'b001
`define 3'b101
LOADBYTEU 3'b011
`define 
LOADHALF 
`define 
LOADHALFU 
`define 
LOADWORD 

