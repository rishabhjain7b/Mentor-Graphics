//Inverter

module inverter
(input a,
 output y);

assign y=~a;
endmodule