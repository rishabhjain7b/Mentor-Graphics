`include"test.sv"

module test1;
test t1;
initial
begin
	t1=new();
	//t1.a=22;
	//t1.b=33;
	t1.display();
end
endmodule
