module multi_array;

//int arr[0:1][0:3]='{2{'{7,3,5,2}}};
int arr[3][4]='{ {2{'{default:7}}} , {1{'{default:5}}} };
initial
begin
	for(int i=0;i<3;i++)
	begin
		for(int j=0;j<4;j++)
		$write("arr[%0d][%0d]=%0d\t",i,j,arr[i][j]);
		$display("");
	end
end
endmodule
