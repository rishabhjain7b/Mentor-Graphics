//buffer
module buffer
(input a,
 output y);

assign y=a;
endmodule