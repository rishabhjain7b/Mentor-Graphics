
`include "alu_packet.sv"
`include "alu_generator.sv"
`include "alu_driver.sv"
`include "alu_intf.sv"
`include "alu_coverage.sv"
`include "alu.sv"
`include "alu_monitor.sv"
`include "alu_scoreboard.sv"
`include "alu_environment.sv"
`include "alu_test.sv"
