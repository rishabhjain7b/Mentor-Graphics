class test;
local int a=2,b;

task display();
begin
	$display("%d %d",a,b);
end
endtask
endclass

