module event_test;
event e1,e2;
initial
begin
	$display("1 before triggered",$time);
	->e1;
	@ e2;
	//wait (e2.triggered);
	$display("1 after triggered",$time);
end
initial
begin
	$display("2 before triggered",$time);
	->e2;
	wait (e1.triggered);
	$display("2 after triggered",$time);
end
endmodule
