// executive preprocessor stage 1

`define CLK_PERIOD 10

`define REGISTER_WIDTH 32
`define INSTR_WIDTH 32
`define IMMEDIATE_WIDTH 16

`define MEM_READ 3'b101
`define MEM_WRITE 3'b100
`define ARITH_LOGIC 3'b001
`define SHIFT_REG 3'b000

// ARITHMETIC 
`define ADD 3'b000
`define HADD 3'b001
`define SUB 3'b010
`define NOT 3'b011
`define AND 3'b100
`define OR 3'b101
`define XOR 3'b110
`define LHG 3'b111
 
// SHIFTING 
`define SHLEFTLOG 3'b000
`define SHLEFTART 3'b001
`define SHRGHTLOG 3'b010
`define SHRGHTART 3'b011
 
// DATA TRANSFER 

`define LOADBYTE 3'b000 
`define LOADBYTEU 3'b100 
`define LOADHALF 3'b001
`define LOADHALFU 3'b101 
`define LOADWORD 3'b011


module preprocessor
(input clock,
 input reset,enable_ex,
 input signed [31:0]src1,src2,imm,mem_data_read_in,
 input [6:0]control_in,
 output mem_data_wr_en,
 output signed [31:0]mem_data_write_out,
 output signed [31:0]aluin1,aluin2,
 output [2:0]operation_out,opselect_out,
 output [4:0]shift_number,
 output enable_arith,enable_shift);
 
 reg signed [31:0]w_aluin1=0;
 reg signed [31:0]w_aluin2=0;
 reg [2:0]w_operation_out=0,w_opselect_out=0;
 reg [4:0]w_shift_number=0;
 reg w_enable_arith=0,w_enable_shift=0;
 
 assign mem_data_write_out=src2,
 	mem_data_wr_en= ((control_in[2:0] == `MEM_WRITE) && (control_in[3] == 1))?1'b1:1'b0;

 assign aluin1=w_aluin1,
 	aluin2=w_aluin2,
 	operation_out=w_operation_out,
 	opselect_out=w_opselect_out,
 	shift_number=w_shift_number,
 	enable_arith=w_enable_arith,
 	enable_shift=w_enable_shift;
 
always @(posedge clock,negedge reset)
begin
	if(!reset)
	begin
		w_aluin1<=0;
		w_aluin2<=0;
		w_operation_out<=0;
		w_opselect_out<=0;
		w_shift_number<=0;
		w_enable_arith<=0;
		w_enable_shift<=0;
	end
	else
	begin
		if(!enable_ex)
		begin
			w_aluin1<=w_aluin1;
			w_aluin2<=w_aluin2;
			w_operation_out<=w_operation_out;
			w_opselect_out<=w_opselect_out;
			w_shift_number<=0;
			w_enable_arith<=0;
			w_enable_shift<=0;
		end
		else
		begin
			w_aluin1<=src1;
			w_operation_out<=control_in[6:4];
			w_opselect_out<=control_in[2:0];
			
			case(control_in[2:0])
			`ARITH_LOGIC:
			begin
				if(control_in[3])
				begin
					w_aluin2<=imm;
					w_shift_number<=0;
					w_enable_arith<=1;
					w_enable_shift<=0;
				end
				
				else
				begin
					w_aluin2<=src2;
					w_shift_number<=0;
					w_enable_arith<=1;
					w_enable_shift<=0;
				end
			end
			
			`MEM_READ:
			begin
				if(control_in[3])
				begin
					w_aluin2<=mem_data_read_in;
					w_shift_number<=0;
					w_enable_arith<=1;
					w_enable_shift<=0;
				end
				
				else
				begin
					w_aluin2<=w_aluin2;
					w_shift_number<=0;
					w_enable_arith<=0;
					w_enable_shift<=0;
				end
			end

			`MEM_WRITE:
			begin
				if(control_in[3])
				begin
					w_aluin2<=w_aluin2;
					w_shift_number<=0;
					w_enable_arith<=0;
					w_enable_shift<=0;
				end
				
				else
				begin
					w_aluin2<=w_aluin2;
					w_shift_number<=0;
					w_enable_arith<=0;
					w_enable_shift<=0;
				end
			end

			`SHIFT_REG:
			begin
				if(control_in[3])
				begin
					w_aluin2<=w_aluin2;
					w_shift_number<=src2[4:0];
					w_enable_arith<=0;
					w_enable_shift<=1;
				end
				
				else
				begin
					w_aluin2<=w_aluin2;
					w_shift_number<=imm[10:6];
					w_enable_arith<=0;
					w_enable_shift<=1;
				end
			end
			endcase
		end
	end
end
endmodule
