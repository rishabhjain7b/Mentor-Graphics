// packet class

class packet;
rand bit [3:0]a,b;
rand bit [2:0]sel;
bit [3:0]s;
bit co;
endclass

