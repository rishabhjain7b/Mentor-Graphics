// packet class

class packet;
rand bit[2:0]a;
rand bit[5:0]b;
endclass

